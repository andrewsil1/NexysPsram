-- +------------------------------------------------------------------------------------------------------------------------------+
-- �                                                   TERMS OF USE: MIT License                                                  �
-- �                                                            																  �
-- +------------------------------------------------------------------------------------------------------------------------------�
-- �Permission is hereby granted, free of charge, to any person obtaining a copy of this software and associated documentation    � 
-- �files (the "Software"), to deal in the Software without restriction, including without limitation the rights to use, copy,    �
-- �modify, merge, publish, distribute, sublicense, and/or sell copies of the Software, and to permit persons to whom the Software�
-- �is furnished to do so, subject to the following conditions:                                                                   �
-- �                                                                                                                              �
-- �The above copyright notice and this permission notice shall be included in all copies or substantial portions of the Software.�
-- �                                                                                                                              �
-- �THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE          �
-- �WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR         �
-- �COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE,   �
-- �ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.                         �
-- +------------------------------------------------------------------------------------------------------------------------------+

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity psram_ip_v1_0_S00_AXI is
	generic (
		-- Users to add parameters here

		-- User parameters ends
		-- Do not modify the parameters beyond this line

		-- Width of ID for for write address, write data, read address and read data
		C_S_AXI_ID_WIDTH	: integer	:= 1;
		-- Width of S_AXI data bus
		C_S_AXI_DATA_WIDTH	: integer	:= 32;
		-- Width of S_AXI address bus
		C_S_AXI_ADDR_WIDTH	: integer	:= 24;
		-- Width of optional user defined signal in write address channel
		C_S_AXI_AWUSER_WIDTH	: integer	:= 0;
		-- Width of optional user defined signal in read address channel
		C_S_AXI_ARUSER_WIDTH	: integer	:= 0;
		-- Width of optional user defined signal in write data channel
		C_S_AXI_WUSER_WIDTH	: integer	:= 0;
		-- Width of optional user defined signal in read data channel
		C_S_AXI_RUSER_WIDTH	: integer	:= 0;
		-- Width of optional user defined signal in write response channel
		C_S_AXI_BUSER_WIDTH	: integer	:= 0
	);
	port (
		-- Users to add ports here

		-- User ports ends
		-- Do not modify the ports beyond this line

		-- Global Clock Signal
		S_AXI_ACLK	: in std_logic;
		-- Global Reset Signal. This Signal is Active LOW
		S_AXI_ARESETN	: in std_logic;
		-- Write Address ID
		S_AXI_AWID	: in std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
		-- Write address
		S_AXI_AWADDR	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
		-- Burst length. The burst length gives the exact number of transfers in a burst
		S_AXI_AWLEN	: in std_logic_vector(7 downto 0);
		-- Burst size. This signal indicates the size of each transfer in the burst
		S_AXI_AWSIZE	: in std_logic_vector(2 downto 0);
		-- Burst type. The burst type and the size information, 
    -- determine how the address for each transfer within the burst is calculated.
		S_AXI_AWBURST	: in std_logic_vector(1 downto 0);
		-- Lock type. Provides additional information about the
    -- atomic characteristics of the transfer.
		S_AXI_AWLOCK	: in std_logic;
		-- Memory type. This signal indicates how transactions
    -- are required to progress through a system.
		S_AXI_AWCACHE	: in std_logic_vector(3 downto 0);
		-- Protection type. This signal indicates the privilege
    -- and security level of the transaction, and whether
    -- the transaction is a data access or an instruction access.
		S_AXI_AWPROT	: in std_logic_vector(2 downto 0);
		-- Quality of Service, QoS identifier sent for each
    -- write transaction.
		S_AXI_AWQOS	: in std_logic_vector(3 downto 0);
		-- Region identifier. Permits a single physical interface
    -- on a slave to be used for multiple logical interfaces.
		S_AXI_AWREGION	: in std_logic_vector(3 downto 0);
		-- Optional User-defined signal in the write address channel.
		S_AXI_AWUSER	: in std_logic_vector(C_S_AXI_AWUSER_WIDTH-1 downto 0);
		-- Write address valid. This signal indicates that
    -- the channel is signaling valid write address and
    -- control information.
		S_AXI_AWVALID	: in std_logic;
		-- Write address ready. This signal indicates that
    -- the slave is ready to accept an address and associated
    -- control signals.
		S_AXI_AWREADY	: out std_logic;
		-- Write Data
		S_AXI_WDATA	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		-- Write strobes. This signal indicates which byte
    -- lanes hold valid data. There is one write strobe
    -- bit for each eight bits of the write data bus.
		S_AXI_WSTRB	: in std_logic_vector((C_S_AXI_DATA_WIDTH/8)-1 downto 0);
		-- Write last. This signal indicates the last transfer
    -- in a write burst.
		S_AXI_WLAST	: in std_logic;
		-- Optional User-defined signal in the write data channel.
		S_AXI_WUSER	: in std_logic_vector(C_S_AXI_WUSER_WIDTH-1 downto 0);
		-- Write valid. This signal indicates that valid write
    -- data and strobes are available.
		S_AXI_WVALID	: in std_logic;
		-- Write ready. This signal indicates that the slave
    -- can accept the write data.
		S_AXI_WREADY	: out std_logic;
		-- Response ID tag. This signal is the ID tag of the
    -- write response.
		S_AXI_BID	: out std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
		-- Write response. This signal indicates the status
    -- of the write transaction.
		S_AXI_BRESP	: out std_logic_vector(1 downto 0);
		-- Optional User-defined signal in the write response channel.
		S_AXI_BUSER	: out std_logic_vector(C_S_AXI_BUSER_WIDTH-1 downto 0);
		-- Write response valid. This signal indicates that the
    -- channel is signaling a valid write response.
		S_AXI_BVALID	: out std_logic;
		-- Response ready. This signal indicates that the master
    -- can accept a write response.
		S_AXI_BREADY	: in std_logic;
		-- Read address ID. This signal is the identification
    -- tag for the read address group of signals.
		S_AXI_ARID	: in std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
		-- Read address. This signal indicates the initial
    -- address of a read burst transaction.
		S_AXI_ARADDR	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
		-- Burst length. The burst length gives the exact number of transfers in a burst
		S_AXI_ARLEN	: in std_logic_vector(7 downto 0);
		-- Burst size. This signal indicates the size of each transfer in the burst
		S_AXI_ARSIZE	: in std_logic_vector(2 downto 0);
		-- Burst type. The burst type and the size information, 
    -- determine how the address for each transfer within the burst is calculated.
		S_AXI_ARBURST	: in std_logic_vector(1 downto 0);
		-- Lock type. Provides additional information about the
    -- atomic characteristics of the transfer.
		S_AXI_ARLOCK	: in std_logic;
		-- Memory type. This signal indicates how transactions
    -- are required to progress through a system.
		S_AXI_ARCACHE	: in std_logic_vector(3 downto 0);
		-- Protection type. This signal indicates the privilege
    -- and security level of the transaction, and whether
    -- the transaction is a data access or an instruction access.
		S_AXI_ARPROT	: in std_logic_vector(2 downto 0);
		-- Quality of Service, QoS identifier sent for each
    -- read transaction.
		S_AXI_ARQOS	: in std_logic_vector(3 downto 0);
		-- Region identifier. Permits a single physical interface
    -- on a slave to be used for multiple logical interfaces.
		S_AXI_ARREGION	: in std_logic_vector(3 downto 0);
		-- Optional User-defined signal in the read address channel.
		S_AXI_ARUSER	: in std_logic_vector(C_S_AXI_ARUSER_WIDTH-1 downto 0);
		-- Write address valid. This signal indicates that
    -- the channel is signaling valid read address and
    -- control information.
		S_AXI_ARVALID	: in std_logic;
		-- Read address ready. This signal indicates that
    -- the slave is ready to accept an address and associated
    -- control signals.
		S_AXI_ARREADY	: out std_logic;
		-- Read ID tag. This signal is the identification tag
    -- for the read data group of signals generated by the slave.
		S_AXI_RID	: out std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
		-- Read Data
		S_AXI_RDATA	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		-- Read response. This signal indicates the status of
    -- the read transfer.
		S_AXI_RRESP	: out std_logic_vector(1 downto 0);
		-- Read last. This signal indicates the last transfer
    -- in a read burst.
		S_AXI_RLAST	: out std_logic;
		-- Optional User-defined signal in the read address channel.
		S_AXI_RUSER	: out std_logic_vector(C_S_AXI_RUSER_WIDTH-1 downto 0);
		-- Read valid. This signal indicates that the channel
    -- is signaling the required read data.
		S_AXI_RVALID	: out std_logic;
		-- Read ready. This signal indicates that the master can
    -- accept the read data and response information.
		S_AXI_RREADY	: in std_logic;
		
    -- Pass physical PSRAM signals up and out		
		MEM_ADDR_OUT  : out std_logic_vector(22 downto 0);  -- To PSRAM address
		MEM_CEN         : out STD_LOGIC;                    -- To PSRAM chip enable
        MEM_OEN         : out STD_LOGIC;                    -- To PSRAM output enable
        MEM_WEN         : out STD_LOGIC;                    -- To PSRAM write enable
        MEM_LBN         : out STD_LOGIC;                    -- To PSRAM low byte write enable
        MEM_UBN         : out STD_LOGIC;                    -- To PSRAM high byte write enable
        MEM_ADV         : out STD_LOGIC;                    -- To PSRAM address valid line
        MEM_CRE         : out STD_LOGIC;
        MEM_DATA_I      : in STD_LOGIC_VECTOR(15 downto 0); -- To PSRAM data bus
        MEM_DATA_O      : out STD_LOGIC_VECTOR(15 downto 0);-- To PSRAM data bus
        MEM_DATA_T      : out STD_LOGIC_VECTOR(15 downto 0)-- To PSRAM data bus
	);
end psram_ip_v1_0_S00_AXI;

architecture arch_imp of psram_ip_v1_0_S00_AXI is

    component AsyncPSRAM is -- Import PSRAM controller module signals
        port(
            sysclk          : in STD_LOGIC;
            rst             : in STD_LOGIC;
            mem_data_wr     : in STD_LOGIC_VECTOR(15 downto 0); 
            mem_addr        : in STD_LOGIC_VECTOR(22 downto 0); 
            mem_byte_en     : in STD_LOGIC_VECTOR(1 downto 0); 
            command         : in STD_LOGIC;                     -- 0 = write, 1 = read
            go              : in STD_LOGIC;                     -- Signals that the command is ready to run.
            mem_idle        : out STD_LOGIC;                    -- 1 = unit is idle, ready for a command, 0 = busy.
            mem_data_rd     : out STD_LOGIC_VECTOR(15 downto 0);-- Contains last read data.
            MEM_ADDR_OUT    : out STD_LOGIC_VECTOR(22 downto 0);-- To PSRAM address bus
            MEM_CEN         : out STD_LOGIC;                    -- To PSRAM chip enable
            MEM_OEN         : out STD_LOGIC;                    -- To PSRAM output enable
            MEM_WEN         : out STD_LOGIC;                    -- To PSRAM write enable
            MEM_LBN         : out STD_LOGIC;                    -- To PSRAM low byte write enable
            MEM_UBN         : out STD_LOGIC;                    -- To PSRAM high byte write enable
            MEM_ADV         : out STD_LOGIC;                    -- To PSRAM address valid line
            MEM_CRE         : out STD_LOGIC;                    -- 
            MEM_DATA_I      : in STD_LOGIC_VECTOR(15 downto 0); -- To PSRAM data bus
            MEM_DATA_O      : out STD_LOGIC_VECTOR(15 downto 0); -- To PSRAM data bus
            MEM_DATA_T      : out STD_LOGIC_VECTOR(15 downto 0) -- To PSRAM data bus
            );
      end component AsyncPSRAM;

	-- AXI4FULL signals
	signal axi_awaddr	: std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
	signal axi_awready	: std_logic;
	signal axi_wready	: std_logic;
	signal axi_bresp	: std_logic_vector(1 downto 0);
	signal axi_buser	: std_logic_vector(C_S_AXI_BUSER_WIDTH-1 downto 0);
	signal axi_bvalid	: std_logic;
	signal axi_araddr	: std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
	signal axi_arready	: std_logic;
	signal axi_rdata	: std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal axi_rresp	: std_logic_vector(1 downto 0);
	signal axi_rlast	: std_logic;
	signal axi_ruser	: std_logic_vector(C_S_AXI_RUSER_WIDTH-1 downto 0);
	signal axi_rvalid	: std_logic;
	-- aw_wrap_en determines wrap boundary and enables wrapping
	signal  aw_wrap_en : std_logic; 
	-- ar_wrap_en determines wrap boundary and enables wrapping
	signal  ar_wrap_en : std_logic;
	-- aw_wrap_size is the size of the write transfer, the
	-- write address wraps to a lower address if upper address
	-- limit is reached
	signal aw_wrap_size : integer;
	-- ar_wrap_size is the size of the read transfer, the
	-- read address wraps to a lower address if upper address
	-- limit is reached
	signal ar_wrap_size : integer;
	-- The axi_awv_awr_flag flag marks the presence of write address valid
	signal axi_awv_awr_flag    : std_logic;
	--The axi_arv_arr_flag flag marks the presence of read address valid
	signal axi_arv_arr_flag    : std_logic;
	-- The axi_awlen_cntr internal write address counter to keep track of beats in a burst transaction
	signal axi_awlen_cntr      : std_logic_vector(7 downto 0);
	signal axi_awlen           : std_logic_vector(7 downto 0); --ANDREWSI added.
	--The axi_arlen_cntr internal read address counter to keep track of beats in a burst transaction
	signal axi_arlen_cntr      : std_logic_vector(7 downto 0);
	signal axi_arlen           : std_logic_vector(7 downto 0); --ANDREWSI added.
	--local parameter for addressing 32 bit / 64 bit C_S_AXI_DATA_WIDTH
	--ADDR_LSB is used for addressing 32/64 bit registers/memories
	--ADDR_LSB = 2 for 32 bits (n downto 2) 
	--ADDR_LSB = 3 for 64 bits (n downto 3)
	constant ADDR_LSB  : integer := (C_S_AXI_DATA_WIDTH/32)+ 1;
	constant OPT_MEM_ADDR_BITS : integer := 7;
	constant low : std_logic_vector (C_S_AXI_ADDR_WIDTH - 1 downto 0) := (others => '0');
	
	------------------------------------------------
    ---- Signals for PSRAM access
    --------------------------------------------------
	signal mem_data_rd, mem_data_wr : std_logic_vector(15 downto 0);
	signal mem_addr : std_logic_vector(22 downto 0);
	signal mem_byte_en : std_logic_vector(1 downto 0);
	signal command, go, mem_idle : std_logic;
	
	------------------------------------------------
	---- Signals for user logic memory space example
	--------------------------------------------------
	signal mem_address : std_logic_vector(22 downto 0);
	signal mem_rden : std_logic;
    signal mem_wren : std_logic;
    
    type state_type is (ST_IDLE, ST_WRITE_L, ST_WRITE_H, ST_READ_L, ST_READ_H);
    signal state, next_state : state_type;
    
begin -- Main Module Code

    -- Instantiate PSRAM controller
    AsyncPSRAMinst : AsyncPSRAM
        port map (
            sysclk => S_AXI_ACLK,
            rst => S_AXI_ARESETN,
            mem_data_wr => mem_data_wr,
            mem_addr => mem_addr,
            mem_byte_en => mem_byte_en,
            command => command,
            go => go,
            mem_idle => mem_idle,
            mem_data_rd => mem_data_rd,
            MEM_ADDR_OUT => MEM_ADDR_OUT,
            MEM_CEN => MEM_CEN,
            MEM_OEN => MEM_OEN,
            MEM_WEN => MEM_WEN,
            MEM_LBN => MEM_LBN,
            MEM_UBN => MEM_UBN,
            MEM_ADV => MEM_ADV,
            MEM_CRE => MEM_CRE,
            MEM_DATA_I => MEM_DATA_I,
            MEM_DATA_O => MEM_DATA_O,
            MEM_DATA_T => MEM_DATA_T
        ); 
	
	-- I/O Connections assignments
	S_AXI_AWREADY <= axi_awready;
	S_AXI_WREADY <= axi_wready;
	S_AXI_BRESP	<= axi_bresp;
	S_AXI_BUSER	<= axi_buser;
	S_AXI_BVALID <= axi_bvalid;
	S_AXI_ARREADY <= axi_arready;
	S_AXI_RDATA	<= axi_rdata;
	S_AXI_RRESP	<= axi_rresp;
	S_AXI_RLAST	<= axi_rlast;
	S_AXI_RUSER	<= axi_ruser;
	S_AXI_RVALID <= axi_rvalid;
	S_AXI_BID <= S_AXI_AWID;
	S_AXI_RID <= S_AXI_ARID;
	aw_wrap_size <= (C_S_AXI_DATA_WIDTH/8 * CONV_INTEGER(S_AXI_AWLEN)); 
	ar_wrap_size <= (C_S_AXI_DATA_WIDTH/8 * CONV_INTEGER(S_AXI_ARLEN)); 
	aw_wrap_en <= '1' when (((axi_awaddr AND CONV_STD_LOGIC_VECTOR(aw_wrap_size,C_S_AXI_ADDR_WIDTH)) XOR CONV_STD_LOGIC_VECTOR(aw_wrap_size,C_S_AXI_ADDR_WIDTH)) = low) else '0';
	ar_wrap_en <= '1' when (((axi_araddr AND CONV_STD_LOGIC_VECTOR(ar_wrap_size,C_S_AXI_ADDR_WIDTH)) XOR CONV_STD_LOGIC_VECTOR(ar_wrap_size,C_S_AXI_ADDR_WIDTH)) = low) else '0';
	S_AXI_BUSER <= (others => '0');

	-- Implement axi_awready generation

	-- axi_awready is asserted for one S_AXI_ACLK clock cycle when both
	-- S_AXI_AWVALID and S_AXI_WVALID are asserted. axi_awready is
	-- de-asserted when reset is low.

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_awready <= '0';
	      axi_awv_awr_flag <= '0';
	    else
	      if (axi_awready = '0' and S_AXI_AWVALID = '1' and axi_awv_awr_flag = '0' and axi_arv_arr_flag = '0') then
	        -- slave is ready to accept an address and
	        -- associated control signals
	        axi_awv_awr_flag  <= '1'; -- used for generation of bresp() and bvalid
	        axi_awready <= '1';
	      elsif (S_AXI_WLAST = '1' and axi_wready = '1') then 
	      -- preparing to accept next address after current write burst tx completion
	        axi_awv_awr_flag  <= '0';
	      else
	        axi_awready <= '0';
	      end if;
	    end if;
	  end if;         
	end process; 
	-- Implement axi_awaddr latching

	-- This process is used to latch the address when both 
	-- S_AXI_AWVALID and S_AXI_WVALID are valid. 

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_awaddr <= (others => '0');
	      axi_awlen_cntr <= (others => '0');
	      axi_awlen <= (others => '0');
	    else
	      if (axi_awready = '0' and S_AXI_AWVALID = '1' and axi_awv_awr_flag = '0') then
	      -- address latching 
	        axi_awaddr <= S_AXI_AWADDR(C_S_AXI_ADDR_WIDTH - 1 downto 0);  ---- start address of transfer
	        axi_awlen_cntr <= (others => '0');
	        axi_awlen <= S_AXI_AWLEN;
	      elsif((axi_awlen_cntr <= axi_awlen) and axi_wready = '1' and S_AXI_WVALID = '1') then     
	        axi_awlen_cntr <= axi_awlen_cntr + '1';

	        case (S_AXI_AWBURST) is
	          when "00" => -- fixed burst
	            -- The write address for all the beats in the transaction are fixed
	            axi_awaddr     <= axi_awaddr;       ----for awsize = 4 bytes (010)
	          when "01" => --incremental burst
	            -- The write address for all the beats in the transaction are increments by awsize
	            axi_awaddr(C_S_AXI_ADDR_WIDTH - 1 downto ADDR_LSB) <= axi_awaddr(C_S_AXI_ADDR_WIDTH - 1 downto ADDR_LSB) + '1';--awaddr aligned to 4 byte boundary
	            axi_awaddr(ADDR_LSB-1 downto 0)  <= (others => '0');  ----for awsize = 4 bytes (010)
	          when "10" => --Wrapping burst
	            -- The write address wraps when the address reaches wrap boundary 
	            if (aw_wrap_en = '1') then
	              axi_awaddr <= axi_awaddr - CONV_STD_LOGIC_VECTOR(aw_wrap_size,C_S_AXI_ADDR_WIDTH);                
	            else 
	              axi_awaddr(C_S_AXI_ADDR_WIDTH - 1 downto ADDR_LSB) <= axi_awaddr(C_S_AXI_ADDR_WIDTH - 1 downto ADDR_LSB) + '1';--awaddr aligned to 4 byte boundary
	              axi_awaddr(ADDR_LSB-1 downto 0)  <= (others => '0');  ----for awsize = 4 bytes (010)
	            end if;
	          when others => --reserved (incremental burst for example)
	            axi_awaddr(C_S_AXI_ADDR_WIDTH - 1 downto ADDR_LSB) <= axi_awaddr(C_S_AXI_ADDR_WIDTH - 1 downto ADDR_LSB) + '1';--for awsize = 4 bytes (010)
	            axi_awaddr(ADDR_LSB-1 downto 0)  <= (others => '0');
	        end case;        
	      end if;
	    end if;
	  end if;
	end process;

	-- Implement write response logic generation

	-- The write response and response valid signals are asserted by the slave 
	-- when axi_wready, S_AXI_WVALID, axi_wready and S_AXI_WVALID are asserted.  
	-- This marks the acceptance of address and indicates the status of 
	-- write transaction.

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_bvalid  <= '0';
	      axi_bresp  <= "00"; --need to work more on the responses
	    else
	      if (axi_awv_awr_flag = '1' and axi_wready = '1' and S_AXI_WVALID = '1' and axi_bvalid = '0' and S_AXI_WLAST = '1' ) then
	        axi_bvalid <= '1';
	        axi_bresp  <= "00"; 
	      elsif (S_AXI_BREADY = '1' and axi_bvalid = '1') then  
	      --check if bready is asserted while bvalid is high)
	        axi_bvalid <= '0';                      
	      end if;
	    end if;
	  end if;         
	end process; 
	-- Implement axi_arready generation

	-- axi_arready is asserted for one S_AXI_ACLK clock cycle when
	-- S_AXI_ARVALID is asserted. axi_awready is 
	-- de-asserted when reset (active low) is asserted. 
	-- The read address is also latched when S_AXI_ARVALID is 
	-- asserted. axi_araddr is reset to zero on reset assertion.

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_arready <= '0';
	      axi_arv_arr_flag <= '0';
	    else
	      if (axi_arready = '0' and S_AXI_ARVALID = '1' and axi_awv_awr_flag = '0' and axi_arv_arr_flag = '0') then
	        axi_arready <= '1';
	        axi_arv_arr_flag <= '1';
	      elsif (axi_rvalid = '1' and S_AXI_RREADY = '1' and (axi_arlen_cntr = axi_arlen)) then 
	      -- preparing to accept next address after current read completion
	        axi_arv_arr_flag <= '0';
	      else
	        axi_arready <= '0';
	      end if;
	    end if;
	  end if;         
	end process; 
	-- Implement axi_araddr latching

	--This process is used to latch the address when both 
	--S_AXI_ARVALID and S_AXI_RVALID are valid. 
	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_araddr <= (others => '0');
	      axi_arlen_cntr <= (others => '0');
	      axi_arlen <= (others => '0');
	      axi_rlast <= '0';
	    else
	      if (axi_arready = '0' and S_AXI_ARVALID = '1' and axi_arv_arr_flag = '0') then
	        -- address latching 
	        axi_araddr <= S_AXI_ARADDR(C_S_AXI_ADDR_WIDTH - 1 downto 0); ---- start address of transfer
	        axi_arlen_cntr <= (others => '0');
	        axi_arlen <= S_AXI_ARLEN;
	        axi_rlast <= '0';
	      elsif((axi_arlen_cntr <= axi_arlen) and axi_rvalid = '1' and S_AXI_RREADY = '1') then     
	        axi_arlen_cntr <= axi_arlen_cntr + '1';
	        axi_rlast <= '0';      
	     
	        case (S_AXI_ARBURST) is
	          when "00" =>  -- fixed burst
	            -- The read address for all the beats in the transaction are fixed
	            axi_araddr     <= axi_araddr;      ----for arsize = 4 bytes (010)
	          when "01" =>  --incremental burst
	            -- The read address for all the beats in the transaction are increments by awsize
	            axi_araddr(C_S_AXI_ADDR_WIDTH - 1 downto ADDR_LSB) <= axi_araddr(C_S_AXI_ADDR_WIDTH - 1 downto ADDR_LSB) + '1'; --araddr aligned to 4 byte boundary
	            axi_araddr(ADDR_LSB-1 downto 0)  <= (others => '0');  ----for awsize = 4 bytes (010)
	          when "10" =>  --Wrapping burst
	            -- The read address wraps when the address reaches wrap boundary 
	            if (ar_wrap_en = '1') then   
	              axi_araddr <= axi_araddr - CONV_STD_LOGIC_VECTOR(ar_wrap_size,C_S_AXI_ADDR_WIDTH);
	            else 
	              axi_araddr(C_S_AXI_ADDR_WIDTH - 1 downto ADDR_LSB) <= axi_araddr(C_S_AXI_ADDR_WIDTH - 1 downto ADDR_LSB) + '1'; --araddr aligned to 4 byte boundary
	              axi_araddr(ADDR_LSB-1 downto 0)  <= (others => '0');  ----for awsize = 4 bytes (010)
	            end if;
	          when others => --reserved (incremental burst for example)
	            axi_araddr(C_S_AXI_ADDR_WIDTH - 1 downto ADDR_LSB) <= axi_araddr(C_S_AXI_ADDR_WIDTH - 1 downto ADDR_LSB) + '1';--for arsize = 4 bytes (010)
			  axi_araddr(ADDR_LSB-1 downto 0)  <= (others => '0');
	        end case;         
	      elsif((axi_arlen_cntr = axi_arlen) and axi_rlast = '0' and axi_arv_arr_flag = '1') then  
	        axi_rlast <= '1';
	      elsif (S_AXI_RREADY = '1') then  
	        axi_rlast <= '0';
	      end if;
	    end if;
	  end if;
	end  process;  
	-- Implement axi_arvalid generation

	-- axi_rvalid is asserted for one S_AXI_ACLK clock cycle when both 
	-- S_AXI_ARVALID and axi_arready are asserted. The slave registers 
	-- data are available on the axi_rdata bus at this instance. The 
	-- assertion of axi_rvalid marks the validity of read data on the 
	-- bus and axi_rresp indicates the status of read transaction.axi_rvalid 
	-- is deasserted on reset (active low). axi_rresp and axi_rdata are 
	-- cleared to zero on reset (active low).  

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then
	    if S_AXI_ARESETN = '0' then
	      axi_rresp  <= "00";
	    else
	      if (axi_arv_arr_flag = '1' and axi_rvalid = '0') then
	        axi_rresp  <= "00"; -- 'OKAY' response
	      end  if;      
	    end if;
	  end if;
	end  process;
	
	-- ------------------------------------------
	-- Code to access PSRAM
	-- ------------------------------------------

    -- Intepret AXI address: LSB is irrelevant since smallest access of PSRAM is 16 bits wide, and unaligned reads need to be realigned first, so
    -- bit 1 is also to be ignored for alignment to 32-bit bus.
  	mem_address <= (axi_araddr(23 downto 2) & '0') when axi_arv_arr_flag = '1' else
	               (axi_awaddr(23 downto 2) & '0') when axi_awv_awr_flag = '1' else
	               (others => '0');
	 
	-- implement PSRAM access wr/rd enable flags based on AXI signals
	  mem_wren <= '1' when (axi_wready = '0' and S_AXI_WVALID = '1' and axi_awv_awr_flag = '1') else '0';
	  mem_rden <= axi_arv_arr_flag;	

   --State-Machine
   MEM_OUTPUT_DECODE: process (S_AXI_ACLK)
   begin
     if (rising_edge(S_AXI_ACLK)) then
       if (S_AXI_ARESETN = '0') then -- RESET
          state <= ST_IDLE;
          axi_wready <= '0';
          axi_rvalid <= '0';
          go <= '0';
          mem_data_wr <= x"0000";
          mem_addr <= (others => '0');
          mem_byte_en <= "00";
          command <= '1';
          axi_rdata <= (others => '0');
       elsif (state = ST_IDLE) then
        state <= next_state;
        axi_wready <= '0';
        axi_rvalid <= '0';
        axi_rdata <= axi_rdata;
        if mem_wren = '1' and S_AXI_WSTRB(1 downto 0) > "00" then -- Go to one of the write states.
            mem_data_wr <= S_AXI_WDATA(15 downto 0);    -- Data for low word
            mem_addr <= mem_address;                    -- Address of 16-bit memory location
            mem_byte_en <= not S_AXI_WSTRB(1 downto 0);   -- Pass on byte write strobes (inverted)
            command <= '0';
            go <= '1';
        elsif mem_wren = '1' and S_AXI_WSTRB(1 downto 0) = "00" then -- In this case the master says not to worry about the lower word, so we can skip it to speed things up.
            mem_data_wr <= S_AXI_WDATA(31 downto 16);    -- Data for high word
            mem_addr <= mem_address + '1';               -- Address of next 16-bit memory location
            mem_byte_en <= not S_AXI_WSTRB(3 downto 2);   -- Pass on byte write strobes (inverted)
            command <= '0';
            go <= '1';
        elsif mem_rden = '1' and axi_rvalid = '0' then -- Perform a read.
            if axi_araddr(1) = '0' then 
               mem_addr <= mem_address;                    
            else -- If bit 1 of the address is high, this is an unaligned read (reading bytes 2 and/or 3), so we don't need to read the low word at all.
               mem_addr <= mem_address + '1';
            end if;            
            mem_data_wr <= (others => '0');
            mem_byte_en <= "00";
            command <= '1';
            go <= '1';
        else
            mem_data_wr <= (others => '0');
            go <= '0';
            mem_addr <= (others => '0');
            mem_byte_en <= "11";
            command <= '1';
        end if;
      elsif (state = ST_WRITE_L) then
        state <= next_state;
        axi_rvalid <= '0';
        go <= '0'; -- Drop go signal after command is acknowledged.
        if mem_idle = '1' then -- Is write complete?
            if S_AXI_WSTRB(3 downto 2) > "00" then
                axi_wready <= '0';                            -- Not done writing yet.
                mem_data_wr <= S_AXI_WDATA(31 downto 16);     -- Data for high word
                mem_addr <= mem_addr + '1';                   -- Address of next 16-bit memory location
                mem_byte_en <= not S_AXI_WSTRB(3 downto 2);   -- Pass on byte write strobes (inverted)
                command <= '0';
                go <= '1';
            else
                axi_wready <= '1'; -- No high word to write, it's complete.
                go <= '0';
                command <= command;
                mem_byte_en <= mem_byte_en;
                mem_addr <= mem_addr;
                mem_data_wr <= mem_data_wr;
            end if;
        end if;       
      elsif (state = ST_WRITE_H) then
        state <= next_state;
        go <= '0';
        axi_rvalid <= '0';
        if mem_idle = '1' and go <= '0' then -- Is write complete?
            axi_wready <= '1';
            mem_data_wr <= (others => '0');
            mem_byte_en <= "11";
            mem_addr <= mem_addr;
            command <= command;
        else
            axi_wready <= axi_wready;
            mem_data_wr <= mem_data_wr;
            mem_byte_en <= mem_byte_en;
            mem_addr <= mem_addr;
            command <= command;
        end if;
      elsif (state = ST_READ_L) then
        state <= next_state;
        axi_rvalid <= '0';
        axi_wready <= '0';
        if mem_idle = '1' then
            axi_rdata(15 downto 0) <= mem_data_rd;
            mem_addr <= mem_addr + '1';
            command <= '1';
            go <= '1';
            mem_data_wr <= (others => '0');
        else
            go <= '0';
            command <= command;
            mem_addr <= mem_addr;
            axi_rdata <= axi_rdata;
            mem_data_wr <= (others => '0');
        end if;
      elsif (state = ST_READ_H) then
         state <= next_state;
         axi_wready <= '0';
         go <= '0';
         if mem_idle = '1' and go = '0' then
            axi_rdata(31 downto 16) <= mem_data_rd;
            axi_rdata(15 downto 0) <= axi_rdata(15 downto 0); -- Keep the prior low word bits!
            axi_rvalid <= '1';
            mem_data_wr <= (others => '0');
            command <= command;
            mem_addr <= mem_addr;
         else
            axi_rdata <= axi_rdata;
            axi_rvalid <= '0';
            mem_data_wr <= (others => '0');
            command <= command;
            mem_addr <= mem_addr;
         end if;
      else -- Invalid state
            state <= ST_IDLE;
            axi_wready <= '0';
            axi_rvalid <= '0';
            go <= '0';
            axi_rdata <= (others => '0');
            mem_data_wr <= (others => '0');
            command <= command;
            mem_addr <= mem_addr;
      end if; 
     end if;
   end process;
 
   NEXT_STATE_DECODE: process (state, mem_wren, mem_rden, mem_idle, go, S_AXI_WSTRB)
   begin
      --declare default state for next_state to avoid latches
      next_state <= state;  --default is to stay in current state
      case (state) is
         when ST_IDLE =>
            if mem_wren = '1' and mem_idle = '0' then -- Wait for PSRAM to acknowledge the operation
                if S_AXI_WSTRB(1 downto 0) > "00" then -- Is there a lower word to write?
                    next_state <= ST_WRITE_L; -- Yes
                else
                    next_state <= ST_WRITE_H; -- No
                end if;
            elsif mem_rden = '1' and mem_idle = '0' then -- Wait for PSRAM to acknowledge the operation
                if axi_araddr(1) = '0' then
                    next_state <= ST_READ_L;  -- Read lower word
                else
                    next_state <= ST_READ_H;  -- Jump straight to reading upper word for 16-bit accesses.
                end if;
            end if;
         when ST_WRITE_L =>
            if mem_idle = '1' then -- Wait for write to complete
                if S_AXI_WSTRB(3 downto 2) > "00" then -- Is there an upper word to write?
                    next_state <= ST_WRITE_H; -- Yes
                else
                    next_state <= ST_IDLE; -- No
                end if;
            end if;
         when ST_WRITE_H => -- Wait for write to complete
            if mem_idle = '1' and go = '0' then -- Wait for write to complete before going on
                next_state <= ST_IDLE;
            end if;
         when ST_READ_L =>
            if mem_idle = '1' then -- Wait for read to complete
                next_state <= ST_READ_H;
            end if;
         when ST_READ_H =>
            if mem_idle = '1' and go = '0' then -- Wait for read to complete before going on
                next_state <= ST_IDLE;
            end if;
      end case;      
   end process;

	-- Add user logic here

	-- User logic ends

end arch_imp;
